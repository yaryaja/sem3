magic
tech scmos
timestamp 1669566722
<< nwell >>
rect -4 57 50 80
rect 89 58 143 82
<< ntransistor >>
rect 10 31 12 42
rect 33 31 35 42
rect 118 29 120 40
<< ptransistor >>
rect 10 63 12 74
rect 33 63 35 74
rect 118 65 120 76
<< ndiffusion >>
rect 3 35 10 42
rect 8 31 10 35
rect 12 31 33 42
rect 35 38 40 42
rect 35 31 44 38
rect 98 35 118 40
rect 98 29 102 35
rect 109 29 118 35
rect 120 34 128 40
rect 135 34 138 40
rect 120 29 138 34
<< pdiffusion >>
rect 9 69 10 74
rect 3 63 10 69
rect 12 70 33 74
rect 12 66 21 70
rect 25 66 33 70
rect 12 63 33 66
rect 35 69 38 74
rect 35 63 44 69
rect 98 71 101 76
rect 107 71 118 76
rect 98 65 118 71
rect 120 72 137 76
rect 120 66 128 72
rect 135 66 137 72
rect 120 65 137 66
<< ndcontact >>
rect 3 31 8 35
rect 40 38 44 42
rect 102 29 109 35
rect 128 34 135 40
<< pdcontact >>
rect 3 69 9 74
rect 21 66 25 70
rect 38 69 44 74
rect 101 71 107 76
rect 128 66 135 72
<< psubstratepcontact >>
rect 10 14 15 18
rect 28 14 32 18
rect 45 14 49 18
rect 61 14 65 18
rect 80 14 84 18
<< nsubstratencontact >>
rect 10 90 15 94
rect 31 90 36 94
rect 54 90 59 94
rect 76 90 80 94
rect 93 90 97 94
<< polysilicon >>
rect 10 74 12 85
rect 33 74 35 85
rect 118 76 120 89
rect 10 42 12 63
rect 33 42 35 63
rect 118 54 120 65
rect 64 49 120 54
rect 118 40 120 49
rect 10 26 12 31
rect 33 26 35 31
rect 118 20 120 29
<< polycontact >>
rect 60 49 64 54
<< metal1 >>
rect 3 90 10 94
rect 15 90 31 94
rect 36 90 54 94
rect 59 90 76 94
rect 80 90 93 94
rect 97 90 108 94
rect 3 74 9 90
rect 38 74 44 90
rect 101 76 107 90
rect 21 54 25 66
rect 128 55 135 66
rect 21 50 60 54
rect 40 49 60 50
rect 128 49 150 55
rect 40 42 44 49
rect 128 40 135 49
rect 3 18 8 31
rect 102 18 108 29
rect 3 14 10 18
rect 15 14 28 18
rect 32 14 45 18
rect 49 14 61 18
rect 65 14 80 18
rect 84 14 108 18
rect 102 12 108 14
<< labels >>
rlabel metal1 22 92 22 92 5 Vdd
rlabel metal1 24 16 24 16 1 Gnd
rlabel polysilicon 10 52 10 52 1 A
rlabel polysilicon 34 47 34 47 1 B
rlabel metal1 48 52 48 52 7 out
rlabel metal1 150 49 150 55 7 output
<< end >>
