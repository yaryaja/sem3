* SPICE3 file created from magicor_gate.ext - technology: scmos


.include 22nm_MGK.pm
.param SUPPLY=1
.param LAMBDA=22n
.param width_N={2*LAMBDA}
.param width_P={2*LAMBDA}
.global gnd vdd 

.option scale=0.01u


v_dd vdd gnd  'SUPPLY'
va A gnd pulse 0 1 0 100p 100p 10n 20n
vb B gnd pulse 0 1 0 100p 100p 20n 40n

M1000 a_n21_45# A Gnd Gnd nmos w=11 l=2
+  ad=231 pd=64 as=77 ps=36
M1001 Vdd B out w_n37_71# pmos w=11 l=2
+  ad=176 pd=76 as=231 ps=64
M1002 out B a_n21_45# Gnd nmos w=11 l=2
+  ad=99 pd=40 as=0 ps=0
M1003 out A Vdd w_n37_71# pmos w=11 l=2
+  ad=0 pd=0 as=0 ps=0
C0 B out 0.24fF
C1 w_n37_71# Vdd 3.38fF
C2 w_n37_71# A 3.18fF
C3 w_n37_71# B 3.18fF
C4 w_n37_71# out 1.13fF



.control
tran 1n 120n
plot  A B+1 out+2
.endc
.end
