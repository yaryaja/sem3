magic
tech scmos
timestamp 1668371028
<< nwell >>
rect -23 11 17 30
rect 23 11 51 29
<< ntransistor >>
rect -11 -10 -9 -4
rect 3 -10 5 -4
rect 37 -10 39 -5
<< ptransistor >>
rect -11 17 -9 23
rect 3 17 5 23
rect 37 17 39 23
<< ndiffusion >>
rect -17 -6 -11 -4
rect -17 -10 -16 -6
rect -12 -10 -11 -6
rect -9 -8 -5 -4
rect -1 -8 3 -4
rect -9 -10 3 -8
rect 5 -6 11 -4
rect 5 -10 6 -6
rect 10 -10 11 -6
rect 23 -6 37 -5
rect 23 -10 28 -6
rect 32 -10 37 -6
rect 39 -9 41 -5
rect 45 -9 51 -5
rect 39 -10 51 -9
<< pdiffusion >>
rect -17 19 -16 23
rect -12 19 -11 23
rect -17 17 -11 19
rect -9 17 3 23
rect 5 21 11 23
rect 5 17 7 21
rect 31 19 32 23
rect 36 19 37 23
rect 31 17 37 19
rect 39 21 45 23
rect 39 17 41 21
<< ndcontact >>
rect -16 -10 -12 -6
rect -5 -8 -1 -4
rect 6 -10 10 -6
rect 28 -10 32 -6
rect 41 -9 45 -5
<< pdcontact >>
rect -16 19 -12 23
rect 7 17 11 21
rect 32 19 36 23
rect 41 17 45 21
<< psubstratepcontact >>
rect -15 -23 -11 -19
rect -7 -23 -3 -19
rect 11 -23 15 -19
rect 21 -23 25 -19
<< nsubstratencontact >>
rect -9 35 -5 39
rect -1 35 3 39
rect 7 35 11 39
rect 19 35 23 39
rect 29 35 33 39
<< polysilicon >>
rect -11 23 -9 31
rect 3 23 5 31
rect 37 23 39 32
rect -11 -4 -9 17
rect 3 -4 5 17
rect 37 9 39 17
rect 25 5 39 9
rect 37 -5 39 5
rect -11 -13 -9 -10
rect 3 -13 5 -10
rect 37 -13 39 -10
<< polycontact >>
rect 21 5 25 9
<< metal1 >>
rect -16 35 -9 39
rect -5 35 -1 39
rect 3 35 7 39
rect 11 35 19 39
rect 23 35 29 39
rect 33 35 36 39
rect -16 23 -12 35
rect 32 23 36 35
rect 7 9 11 17
rect 7 8 21 9
rect -5 5 21 8
rect 41 5 45 17
rect -5 -4 -1 5
rect 41 1 55 5
rect 41 -5 45 1
rect -16 -19 -12 -10
rect 6 -19 10 -10
rect 28 -19 32 -10
rect -20 -23 -15 -19
rect -11 -23 -7 -19
rect -3 -23 11 -19
rect 15 -23 21 -19
rect 25 -23 32 -19
<< labels >>
rlabel metal1 -1 -21 -1 -21 1 GND
rlabel metal1 -15 37 -15 37 5 VDD
rlabel polysilicon -10 8 -10 8 1 A
rlabel polysilicon 4 9 4 9 1 B
rlabel metal1 52 3 52 3 7 output
<< end >>
