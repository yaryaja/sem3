magic
tech scmos
timestamp 1668121591
<< metal1 >>
rect -17 102 0 106
rect -46 14 -39 19
rect -17 9 -12 102
rect 114 99 137 103
rect -46 4 -12 9
rect -17 -52 -12 4
rect -7 29 0 33
rect -7 19 -3 29
rect -7 -45 -3 14
rect 117 2 137 6
rect -7 -49 42 -45
rect -17 -56 42 -52
rect 117 -55 121 2
rect 107 -59 121 -55
<< metal2 >>
rect -34 14 -7 19
<< m2contact >>
rect -39 14 -34 19
rect -7 14 -3 19
use XOR  XOR_0
timestamp 1668121591
transform 1 0 15 0 1 92
box -15 -92 99 77
use AND  AND_0
timestamp 1668121591
transform 1 0 41 0 1 -86
box 0 0 66 83
<< end >>
