TEST MULTIPLIER
***SETUP***
.INCLUDE TSMC_180nm.txt
.INCLUDE multiplier.sub
.PARAM SUPPLY = 1
.PARAM LAMBDA = 0.18u
.PARAM width_N = {12*LAMBDA}
.PARAM width_P = {2*width_N}
.GLOBAL GND VDD

VDS VDD GND 'SUPPLY'

X1 A0 A1 A2 A3 B0 B1 B2 B3 P0 P1 P2 P3 P4 P5 P6 P7 VDD GND multi_mag

***INPUT***
VA0 A0 GND PULSE(0 1 0 100p 100p 10n 20n)
VA1 A1 GND PULSE(0 1 0 100p 100p 10n 20n)
VA2 A2 GND PULSE(0 1 0 100p 100p 10n 20n)
VA3 A3 GND PULSE(0 1 0 100p 100p 10n 20n)
VB0 B0 GND PULSE(0 1 0 100p 100p 20n 40n)
VB1 B1 GND PULSE(0 1 0 100p 100p 20n 40n)
VB2 B2 GND PULSE(0 1 0 100p 100p 20n 40n)
VB3 B3 GND PULSE(0 1 0 100p 100p 20n 40n)

.TRAN 100p 40n

***ANALYSIS***
.CONTROL
	run
	plot v(P0) v(P1)+2 v(P2)+4 v(P3)+6 v(P4)+8 v(P5)+10 v(P6)+12 v(P7)+14
.ENDC

.END
