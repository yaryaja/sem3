magic
tech scmos
timestamp 1669340375
<< nwell >>
rect 0 0 32 32
<< polysilicon >>
rect 11 26 13 29
rect 19 26 21 29
rect 11 -9 13 6
rect 11 -23 13 -13
rect 19 -16 21 6
rect 19 -23 21 -20
rect 11 -46 13 -43
rect 19 -46 21 -43
<< ndiffusion >>
rect 10 -43 11 -23
rect 13 -43 19 -23
rect 21 -43 24 -23
<< pdiffusion >>
rect 10 6 11 26
rect 13 6 14 26
rect 18 6 19 26
rect 21 6 22 26
<< metal1 >>
rect 0 30 32 33
rect 6 26 10 30
rect 22 26 26 30
rect 14 -2 18 6
rect 14 -6 32 -2
rect -1 -13 9 -9
rect -1 -20 17 -16
rect 24 -19 32 -6
rect 24 -23 28 -19
rect 6 -47 10 -43
rect -1 -50 32 -47
<< ntransistor >>
rect 11 -43 13 -23
rect 19 -43 21 -23
<< ptransistor >>
rect 11 6 13 26
rect 19 6 21 26
<< polycontact >>
rect 9 -13 13 -9
rect 17 -20 21 -16
<< ndcontact >>
rect 6 -43 10 -23
rect 24 -43 28 -23
<< pdcontact >>
rect 6 6 10 26
rect 14 6 18 26
rect 22 6 26 26
<< labels >>
rlabel metal1 13 32 22 33 5 vdd
rlabel metal1 10 -49 19 -48 1 gnd
<< end >>
